`define NVDLA_MAC_ATOMIC_C_SIZE 8
`define NVDLA_MAC_ATOMIC_K_SIZE 8
`define NVDLA_MEMORY_ATOMIC_SIZE 32
`define NVDLA_MAX_BATCH_SIZE 32
`define NVDLA_CBUF_BANK_NUMBER 16
`define NVDLA_CBUF_BANK_WIDTH 64
`define NVDLA_CBUF_BANK_DEPTH 512
`define NVDLA_SDP_BS_THROUGHPUT 1
`define NVDLA_SDP_BN_THROUGHPUT 1
`define NVDLA_SDP_EW_THROUGHPUT 4
`define NVDLA_PDP_THROUGHPUT 1
`define NVDLA_CDP_THROUGHPUT 1
`define NVDLA_PRIMARY_MEMIF_LATENCY 1200
`define NVDLA_SECONDARY_MEMIF_LATENCY 128
`define NVDLA_PRIMARY_MEMIF_MAX_BURST_LENGTH 1
`define NVDLA_PRIMARY_MEMIF_WIDTH 512
`define NVDLA_SECONDARY_MEMIF_MAX_BURST_LENGTH 4
`define NVDLA_SECONDARY_MEMIF_WIDTH 512
